* C:\Users\Vivobook\AppData\Roaming\SPB_Data\eSim-Workspace\Multiplexer\Multiplexer.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 03/03/22 14:55:17

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U3  Net-_U3-Pad1_ Net-_U3-Pad2_ Net-_U3-Pad3_ Net-_U3-Pad4_ sensoham_2to1mux		
U5  i0 i1 sel Net-_U3-Pad1_ Net-_U3-Pad2_ Net-_U3-Pad3_ adc_bridge_3		
U6  Net-_U3-Pad4_ Y dac_bridge_1		
v1  i0 GND pulse		
v2  i1 GND pulse		
v3  sel GND pulse		
R1  Y GND 1k		
U1  i0 plot_v1		
U2  i1 plot_v1		
U4  sel plot_v1		
U7  ? plot_v1		

.end
